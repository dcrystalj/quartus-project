library verilog;
use verilog.vl_types.all;
entity trifid_vlg_vec_tst is
end trifid_vlg_vec_tst;
