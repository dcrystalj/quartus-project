module test3_a(q, a);
output [15:0] q;
input [7:0] a;

assign q = a * 215;

endmodule