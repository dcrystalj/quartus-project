module test3_c(q, a);
output [15:0] q;
input [7:0] a;

assign q = a * 64;

endmodule