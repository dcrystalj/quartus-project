module mod


endmodule